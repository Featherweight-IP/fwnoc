
/****************************************************************************
 * fwnoc_router_arb.v
 ****************************************************************************/

  
/**
 * Module: fwnoc_router_arb
 * 
 * TODO: Add module documentation
 */
module fwnoc_router_arb;


endmodule


