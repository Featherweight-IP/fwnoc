
/****************************************************************************
 * fwnoc.v
 ****************************************************************************/

  
/**
 * Module: fwnoc
 * 
 * TODO: Add module documentation
 */
module fwnoc #(
		parameter X_SIZE=2,
		parameter Y_SIZE=1,
		) (
		);


endmodule


